-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Tuesday, September 11, 2012 16:13:27 Pakistan Standard Time

